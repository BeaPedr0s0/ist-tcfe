.OP
R1 1 2 1.041113e+03 
R2 3 2 2.099452e+03 
R3 2 5 3.131091e+03 
R4 5 0 4.119470e+03 
R5 5 6 3.115588e+03 
R6 9 7 2.047994e+03 
R7 7 8 1.027544e+03 
Vs 1 0 5.068716e+00 
Ve 0 9 0V 
Hd 5 8 Ve 8.115684e+03 
Gb 6 3 (2,5) 7.287471e-03 
.END

