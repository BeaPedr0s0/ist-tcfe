.OP

*INDEPENDENT VOLTAGE SOURCE, CONNECTED TO GROUND. AND NODE X. VALUE IN VOLTS.
Vs 1 0 5.068716e+00 

*RESISTORS, CONNECTED BETWEEN THE NODES X X. RESISTANCE VALUE IN OHM.
R1 1 2 1.041113e+03 
R2 3 2 2.099452e+03 
R3 2 5 3.131091e+03 
R4 5 0 4.119470e+03 
R5 5 6 3.115588e+03 
R6 9 0 2.047994e+03 
R7 7 8 1.027544e+03 

*DEPENDENT CURRENT SOURCE. CONNECTED TO NODES X & X. DEPENDS OF THE VOLTAGE BETWEEN THE NODES 1 AND 4. VALUE AMPLIFIED BY CONSTANT Z. VALUE IN AMPERES.
Gb 6 3 (2,5) 7.287471e-03 

*DEPENDENT VOLTAGE SOURCE. CONNECTED TO NODES X & X . DEPENDS OF THE CURRENT THATS FLOWS IN THE VAUX SOURCE. IS AMPLIFIED BY CONSTANTE Y. VALUE IN VOLTS.
Hd 5 8 Vaux 8.115684e+03 

*INDEPENDENT VOLTAGE SOURCE TO USE IN THE DEPENDENT VOLTAGE SOURCE. CONNECTED TO NODES X & X. VALUE = 0 VOLTS
Vaux 9 7 0 

*CAPACITOR. CONNECTED TO NODES X & X. VALUE = 0 VOLTS
C1 6 8 1.041275e-06 

.END

