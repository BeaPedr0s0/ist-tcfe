.OP

Vcc vcc 0 12 
Vin in 0 0 ac 1.0 sin(0 10m 1k) 
R_in in in2 100

*input  coupling capacitor
C_i in2 base 1.9u 

*bias circuit
R_1 vcc base 76000 
R_2 base 0 19000 

*gain stage
Q1 coll base emit BC547A
R_c vcc coll 20000
R_e emit 0 3900

*bypass capacitor
C_b emit 0 1u

*output stage
Q2 0 coll emit2 BC557A
R_out emit2 vcc 100

*output coupling capacitor
C_out emit2 out 1u

*load
R_L out 0 8

.END

