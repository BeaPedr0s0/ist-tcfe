*
* NGSPICE simulation script lab1
* Group 28
*


.options savecurrents

* supply voltage
Vcc vcc 0 10.0

* input voltage source
Va 0 3 5.06871572779
R1 1 0 1.04111259479k
R2 2 1 2.09945227782k
R3 1 4 3.13109125645k
R4 3 4 4.11947040212k
R5 4 5 3.1155879392k
R6 3 8 2.04799381798k
R7 6 7 1.02754401839k
Id 7 5 1.04127523824m
Gb 5 2 (1,4) 7.28747116393m
Hc 4 7 Vb 8.11568444746m
Vb 8 6  0

.model group 28

.control

op

echo "********************************************"
echo  "Operating point"
echo "********************************************"

echo  "op_TAB"
print all
echo  "op_END"

.endc

.end

