.OP

Vcc vcc 0 12
Vin in 0 0 
Rin in in2 100 

*input  coupling capacitor
Ci in2 base 1.9u 

*bias circuit
R1 vcc base 76000 
R2 base 0 19000 

*gain stage
Q1 coll base emit BC547A
Rc vcc coll 20000
Re emit 0 3900

*bypass capacitor
Cb emit 0 1.0u

*output stage
Q2 0 coll emit2 BC557A
Rout emit2 vcc 100

*output coupling capacitor
Co emit2 out 1u

*fonte de teste
VL out 0 ac 1.0 sin(0 10m 1k)

.END

